-- FSM
