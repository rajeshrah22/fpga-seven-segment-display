-- This is the toplevel
