-- Display FSM
