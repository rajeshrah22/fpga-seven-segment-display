-- FSM

