-- seven segment driver
